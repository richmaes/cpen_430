`define USE_ASYNC_RST
